CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
250 220 30 140 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 438 253 0 1 11
0 6
0
0 0 21104 270
2 0V
-6 -16 8 -8
2 I0
-6 -21 8 -13
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7574 0 0
2
5.89787e-315 5.36716e-315
0
13 Logic Switch~
5 528 252 0 1 11
0 5
0
0 0 21104 270
2 0V
-6 -16 8 -8
2 I1
-6 -21 8 -13
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
881 0 0
2
5.89787e-315 5.3568e-315
0
13 Logic Switch~
5 264 425 0 1 11
0 9
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 A0
-6 -16 8 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
361 0 0
2
5.89787e-315 5.34643e-315
0
13 Logic Switch~
5 265 504 0 1 11
0 19
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 CS
-6 -16 8 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8203 0 0
2
5.89787e-315 5.32571e-315
0
13 Logic Switch~
5 265 529 0 1 11
0 18
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 RD
-6 -16 8 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8173 0 0
2
5.89787e-315 5.30499e-315
0
13 Logic Switch~
5 265 554 0 1 11
0 17
0
0 0 21104 0
2 0V
-6 -16 8 -8
2 OE
-6 -16 8 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3731 0 0
2
5.89787e-315 5.26354e-315
0
13 Logic Switch~
5 635 250 0 1 11
0 7
0
0 0 21104 270
2 0V
-6 -16 8 -8
2 I2
-6 -21 8 -13
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
938 0 0
2
5.89787e-315 0
0
8 2-In OR~
219 498 516 0 3 22
0 30 31 13
0
0 0 112 270
6 74LS32
-21 -24 21 -16
2 A3
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
7731 0 0
2
5.89787e-315 5.47207e-315
0
12 D Flip-Flop~
219 466 327 0 4 9
0 6 4 33 32
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3808 0 0
2
5.89787e-315 5.47077e-315
0
9 3-In AND~
219 384 639 0 4 22
0 18 19 17 16
0
0 0 624 0
5 74F11
-18 -28 17 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 5 0
1 U
8679 0 0
2
5.89787e-315 5.46818e-315
0
9 2-In AND~
219 348 446 0 3 22
0 19 20 8
0
0 0 112 90
5 74F08
-18 -24 17 -16
4 BITD
-15 -34 13 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
3693 0 0
2
5.89787e-315 5.46559e-315
0
9 Inverter~
13 353 486 0 2 22
0 18 20
0
0 0 112 90
5 74F04
-18 -19 17 -11
3 U7C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 7 0
1 U
3922 0 0
2
5.89787e-315 5.463e-315
0
9 Inverter~
13 324 354 0 2 22
0 9 3
0
0 0 112 90
5 74F04
-18 -19 17 -11
3 U7D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 7 0
1 U
3897 0 0
2
5.89787e-315 5.46041e-315
0
12 D Flip-Flop~
219 467 425 0 4 9
0 6 2 34 29
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U9
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3422 0 0
2
5.89787e-315 5.45782e-315
0
9 2-In AND~
219 393 407 0 3 22
0 8 9 2
0
0 0 112 0
5 74F08
-18 -24 17 -16
5 BIT2A
-18 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
8941 0 0
2
5.89787e-315 5.45523e-315
0
12 D Flip-Flop~
219 566 326 0 4 9
0 5 4 35 28
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3861 0 0
2
5.89787e-315 5.45264e-315
0
12 D Flip-Flop~
219 567 427 0 4 9
0 5 2 36 25
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U8
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
930 0 0
2
5.89787e-315 5.45005e-315
0
9 2-In AND~
219 512 370 0 3 22
0 32 3 30
0
0 0 112 270
5 74F08
-18 -24 17 -16
5 BIT3A
-18 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
5194 0 0
2
5.89787e-315 5.44746e-315
0
9 2-In AND~
219 494 480 0 3 22
0 29 9 31
0
0 0 112 270
5 74F08
-18 -24 17 -16
5 BIT3B
-18 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
9343 0 0
2
5.89787e-315 5.44487e-315
0
9 2-In AND~
219 620 370 0 3 22
0 28 3 27
0
0 0 112 270
5 74F08
-18 -24 17 -16
5 BIT3C
-18 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
5701 0 0
2
5.89787e-315 5.44228e-315
0
8 2-In OR~
219 606 516 0 3 22
0 27 26 14
0
0 0 112 270
6 74LS32
-21 -24 21 -16
2 A2
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
6934 0 0
2
5.89787e-315 5.43969e-315
0
9 2-In AND~
219 602 480 0 3 22
0 25 9 26
0
0 0 112 270
5 74F08
-18 -24 17 -16
5 BIT3D
-18 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
5845 0 0
2
5.89787e-315 5.4371e-315
0
12 D Flip-Flop~
219 668 326 0 4 9
0 7 4 37 24
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9508 0 0
2
5.89787e-315 5.43451e-315
0
12 D Flip-Flop~
219 669 426 0 4 9
0 7 2 38 21
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6986 0 0
2
5.89787e-315 5.43192e-315
0
8 2-In OR~
219 716 516 0 3 22
0 23 22 15
0
0 0 112 270
6 74LS32
-21 -24 21 -16
2 A1
-7 -34 7 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
8935 0 0
2
5.89787e-315 5.42933e-315
0
9 2-In AND~
219 730 365 0 3 22
0 24 3 23
0
0 0 112 270
5 74F08
-18 -24 17 -16
5 BIT4A
-18 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
329 0 0
2
5.89787e-315 5.42414e-315
0
9 2-In AND~
219 712 481 0 3 22
0 21 9 22
0
0 0 112 270
5 74F08
-18 -24 17 -16
5 BIT4B
-18 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
7213 0 0
2
5.89787e-315 5.41896e-315
0
14 Logic Display~
6 858 550 0 1 2
10 11
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 D2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8696 0 0
2
5.89787e-315 5.41378e-315
0
14 Logic Display~
6 858 583 0 1 2
10 12
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 D1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3912 0 0
2
5.89787e-315 5.4086e-315
0
14 Logic Display~
6 858 616 0 1 2
10 10
0
0 0 53856 270
6 100MEG
3 -16 45 -8
2 D0
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3882 0 0
2
5.89787e-315 5.40342e-315
0
10 Buffer 3S~
219 783 554 0 3 22
0 15 16 11
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
4408 0 0
2
5.89787e-315 5.39824e-315
0
10 Buffer 3S~
219 782 587 0 3 22
0 14 16 12
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
9377 0 0
2
5.89787e-315 5.39306e-315
0
10 Buffer 3S~
219 782 620 0 3 22
0 13 16 10
0
0 0 112 0
8 BUFFER3S
-27 -51 29 -43
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 9 10 8 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
4560 0 0
2
5.89787e-315 5.38788e-315
0
9 2-In AND~
219 391 309 0 3 22
0 3 8 4
0
0 0 112 0
5 74F08
-18 -24 17 -16
5 BIT4C
-18 -34 17 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
6816 0 0
2
5.89787e-315 5.37752e-315
0
50
0 0 2 0 0 4224 0 0 0 2 17 3
536 436
439 436
439 407
2 2 2 0 0 0 0 24 17 0 0 6
645 408
626 408
626 436
536 436
536 409
543 409
2 0 3 0 0 4096 0 18 0 0 5 2
501 348
501 336
2 0 3 0 0 0 0 20 0 0 5 2
609 348
609 336
2 2 3 0 0 4224 0 13 26 0 0 3
327 336
719 336
719 343
0 2 4 0 0 4096 0 0 23 7 0 4
536 331
639 331
639 308
644 308
0 2 4 0 0 8320 0 0 16 8 0 5
424 309
424 331
536 331
536 308
542 308
2 3 4 0 0 0 0 9 34 0 0 2
442 309
412 309
1 0 5 0 0 4096 0 16 0 0 49 2
542 290
527 290
1 0 6 0 0 4096 0 9 0 0 50 2
442 291
438 291
1 0 7 0 0 4096 0 23 0 0 39 4
644 290
639 290
639 289
635 289
2 1 3 0 0 0 0 13 34 0 0 3
327 336
327 300
367 300
0 2 8 0 0 4224 0 0 34 14 0 3
347 397
347 318
367 318
1 3 8 0 0 0 0 15 11 0 0 5
369 398
347 398
347 397
347 397
347 422
0 0 9 0 0 8320 0 0 0 16 41 3
365 416
365 445
483 445
0 2 9 0 0 0 0 0 15 33 0 2
327 416
369 416
3 2 2 0 0 0 0 15 14 0 0 2
414 407
443 407
3 1 10 0 0 4224 0 33 30 0 0 2
797 620
842 620
1 3 11 0 0 4224 0 28 31 0 0 2
842 554
798 554
3 1 12 0 0 4224 0 32 29 0 0 2
797 587
842 587
1 3 13 0 0 4224 0 33 8 0 0 3
767 620
501 620
501 546
3 1 14 0 0 8320 0 21 32 0 0 3
609 546
609 587
767 587
3 1 15 0 0 8320 0 25 31 0 0 3
719 546
719 554
768 554
0 2 16 0 0 4096 0 0 31 25 0 3
807 603
807 565
783 565
0 2 16 0 0 0 0 0 32 26 0 5
782 639
807 639
807 601
782 601
782 598
4 2 16 0 0 4224 0 10 33 0 0 3
405 639
782 639
782 631
1 3 17 0 0 8320 0 6 10 0 0 4
277 554
332 554
332 648
360 648
0 1 18 0 0 4224 0 0 10 30 0 3
355 529
355 630
360 630
0 2 19 0 0 4224 0 0 10 31 0 3
338 504
338 639
360 639
1 1 18 0 0 0 0 5 12 0 0 3
277 529
356 529
356 504
1 1 19 0 0 0 0 4 11 0 0 3
277 504
338 504
338 467
2 2 20 0 0 4224 0 12 11 0 0 2
356 468
356 467
1 1 9 0 0 0 0 13 3 0 0 3
327 372
327 425
276 425
0 2 9 0 0 0 0 0 27 41 0 4
591 445
591 444
701 444
701 459
4 1 21 0 0 8320 0 24 27 0 0 3
693 390
719 390
719 459
3 2 22 0 0 4224 0 27 25 0 0 2
710 504
710 500
3 1 23 0 0 4224 0 26 25 0 0 2
728 388
728 500
1 4 24 0 0 4224 0 26 23 0 0 3
737 343
737 290
692 290
1 1 7 0 0 4224 0 7 24 0 0 3
635 262
635 390
645 390
1 4 25 0 0 4224 0 22 17 0 0 3
609 458
609 391
591 391
2 2 9 0 0 0 0 22 19 0 0 4
591 458
591 445
483 445
483 458
3 2 26 0 0 4224 0 22 21 0 0 2
600 503
600 500
1 3 27 0 0 4224 0 21 20 0 0 2
618 500
618 393
4 1 28 0 0 8320 0 16 20 0 0 3
590 290
627 290
627 348
4 1 29 0 0 8320 0 14 19 0 0 3
491 389
501 389
501 458
3 1 30 0 0 4224 0 18 8 0 0 2
510 393
510 500
2 3 31 0 0 4224 0 8 19 0 0 2
492 500
492 503
4 1 32 0 0 8320 0 9 18 0 0 3
490 291
519 291
519 348
1 1 5 0 0 12416 0 2 17 0 0 5
528 264
528 290
527 290
527 391
543 391
1 1 6 0 0 4224 0 1 14 0 0 3
438 265
438 389
443 389
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
