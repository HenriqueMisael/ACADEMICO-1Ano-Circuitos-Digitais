CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1155 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
48 C:\Program Files\CircuitMaker 2000 Trial\BOM.DAT
0 7
3 3 0.500000 0.168350
1164 80 1364 747
9437202 0
0
6 Title:
5 Name:
0
0
0
42
10 2-In XNOR~
219 735 185 0 3 22
0 7 10 25
0
0 0 96 270
4 4077
-7 -24 21 -16
4 U11A
30 -9 58 -1
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
5652 0 0
2
42737.8 41
0
5 4030~
219 695 181 0 3 22
0 7 10 26
0
0 0 96 270
4 4030
-7 -24 21 -16
4 U10A
27 -6 55 2
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
4925 0 0
2
42737.8 40
0
9 2-In NOR~
219 652 181 0 3 22
0 7 10 27
0
0 0 96 270
4 7428
-14 -24 14 -16
3 U8A
31 -10 52 -2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
8917 0 0
2
42737.8 39
0
8 2-In OR~
219 604 181 0 3 22
0 7 10 28
0
0 0 96 270
5 74F32
-18 -24 17 -16
3 U1C
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
387 0 0
2
42737.8 38
0
9 2-In AND~
219 484 184 0 3 22
0 7 10 30
0
0 0 96 270
5 74F08
-18 -24 17 -16
2 A5
-8 -34 6 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3329 0 0
2
42737.8 37
0
5 4011~
219 532 186 0 3 22
0 7 10 29
0
0 0 96 270
4 4011
-7 -24 21 -16
3 U9A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 10 0
1 U
515 0 0
2
42737.8 36
0
9 Inverter~
13 847 331 0 2 22
0 23 24
0
0 0 96 180
6 74LS04
-21 -19 21 -11
2 A4
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
7502 0 0
2
42737.8 35
0
9 Inverter~
13 847 368 0 2 22
0 21 22
0
0 0 96 180
6 74LS04
-21 -19 21 -11
2 A3
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
8483 0 0
2
42737.8 34
0
9 Inverter~
13 847 410 0 2 22
0 2 12
0
0 0 96 180
6 74LS04
-21 -19 21 -11
2 A2
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
3730 0 0
2
42737.8 33
0
5 4082~
219 452 475 0 5 22
0 2 22 24 11 39
0
0 0 96 270
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
7176 0 0
2
42737.8 32
0
5 4082~
219 408 475 0 5 22
0 12 22 24 11 40
0
0 0 96 270
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
3493 0 0
2
42737.8 31
0
5 4082~
219 498 476 0 5 22
0 12 21 24 30 38
0
0 0 96 270
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
9394 0 0
2
42737.8 30
0
5 4082~
219 540 476 0 5 22
0 2 21 29 24 37
0
0 0 96 270
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
9594 0 0
2
42737.8 29
0
5 4082~
219 604 476 0 5 22
0 12 28 22 23 36
0
0 0 96 270
4 4082
-7 -24 21 -16
3 U7A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
8880 0 0
2
42737.8 28
0
5 4082~
219 647 476 0 5 22
0 27 2 22 23 35
0
0 0 96 270
4 4082
-7 -24 21 -16
3 U7B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
3776 0 0
2
42737.8 27
0
5 4082~
219 686 476 0 5 22
0 26 12 21 23 34
0
0 0 96 270
4 4082
-7 -24 21 -16
4 U12A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
6204 0 0
2
42737.8 26
0
5 4082~
219 730 476 0 5 22
0 25 2 21 23 33
0
0 0 96 270
4 4082
-7 -24 21 -16
4 U12B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 13 0
1 U
5109 0 0
2
42737.8 25
0
14 Logic Display~
6 497 587 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 S
-3 -21 4 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7406 0 0
2
42737.8 24
0
8 2-In OR~
219 550 592 0 3 22
0 32 31 41
0
0 0 96 270
5 74F32
-18 -24 17 -16
3 U1D
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9403 0 0
2
42737.8 23
0
8 4-In OR~
219 467 533 0 5 22
0 37 38 39 40 31
0
0 0 96 270
4 4072
-14 -24 14 -16
3 U6A
26 -5 47 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 14 0
1 U
3169 0 0
2
42737.8 22
0
8 4-In OR~
219 664 539 0 5 22
0 33 34 35 36 32
0
0 0 96 270
4 4072
-14 -24 14 -16
3 U6B
26 -5 47 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 14 0
1 U
7554 0 0
2
42737.8 21
0
5 4030~
219 290 143 0 3 22
0 7 10 20
0
0 0 96 270
4 4030
-7 -24 21 -16
4 U10B
27 -6 55 2
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
5587 0 0
2
42737.8 20
0
5 4030~
219 281 187 0 3 22
0 20 8 11
0
0 0 96 270
4 4030
-7 -24 21 -16
4 U10C
27 -6 55 2
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 11 0
1 U
7462 0 0
2
42737.8 19
0
9 2-In AND~
219 255 144 0 3 22
0 7 8 18
0
0 0 96 270
5 74F08
-18 -24 17 -16
3 A1A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
8620 0 0
2
42737.8 18
0
9 2-In AND~
219 223 144 0 3 22
0 10 8 19
0
0 0 96 270
5 74F08
-18 -24 17 -16
3 A1B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
5427 0 0
2
42737.8 17
0
9 2-In AND~
219 337 144 0 3 22
0 7 10 17
0
0 0 96 270
5 74F08
-18 -24 17 -16
3 A1C
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
4883 0 0
2
42737.8 16
0
8 3-In OR~
219 250 235 0 4 22
0 17 18 19 13
0
0 0 96 270
4 4075
-14 -24 14 -16
3 U2A
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 7 0
1 U
5670 0 0
2
42737.8 15
0
14 Logic Display~
6 469 587 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
4 Cout
-13 -21 15 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5880 0 0
2
42737.8 14
0
8 2-In OR~
219 416 612 0 3 22
0 15 14 16
0
0 0 96 0
5 74F32
-18 -24 17 -16
3 U5A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
4285 0 0
2
42737.8 13
0
9 2-In AND~
219 264 456 0 3 22
0 12 13 15
0
0 0 96 270
5 74F08
-18 -24 17 -16
3 A1D
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3931 0 0
2
42737.8 12
0
9 2-In AND~
219 230 621 0 3 22
0 2 3 14
0
0 0 96 0
5 74F08
-18 -24 17 -16
3 A6A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
858 0 0
2
42737.8 11
0
9 2-In AND~
219 169 217 0 3 22
0 7 8 4
0
0 0 96 270
5 74F08
-18 -24 17 -16
3 A6D
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
4671 0 0
2
42737.8 10
0
9 2-In AND~
219 135 218 0 3 22
0 7 9 5
0
0 0 96 270
5 74F08
-18 -24 17 -16
3 A6C
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
674 0 0
2
42737.8 9
0
9 2-In AND~
219 101 218 0 3 22
0 9 8 6
0
0 0 96 270
5 74F08
-18 -24 17 -16
3 A6B
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
3611 0 0
2
42737.8 8
0
9 Inverter~
13 173 65 0 2 22
0 10 9
0
0 0 96 180
6 74LS04
-21 -19 21 -11
2 AF
-7 -29 7 -21
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
8345 0 0
2
42737.8 7
0
8 3-In OR~
219 130 285 0 4 22
0 4 5 6 3
0
0 0 96 270
4 4075
-14 -24 14 -16
3 U2B
28 -7 49 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 7 0
1 U
7818 0 0
2
42737.8 6
0
13 Logic Switch~
5 368 30 0 1 11
0 7
0
0 0 21216 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8365 0 0
2
42737.8 5
0
13 Logic Switch~
5 331 32 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21216 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6800 0 0
2
42737.8 4
0
13 Logic Switch~
5 898 307 0 1 11
0 23
0
0 0 21216 180
2 0V
-6 -16 8 -8
2 F0
-6 -16 8 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4638 0 0
2
42737.8 3
0
13 Logic Switch~
5 898 344 0 1 11
0 21
0
0 0 21216 180
2 0V
-6 -16 8 -8
2 F1
-6 -16 8 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8465 0 0
2
42737.8 2
0
13 Logic Switch~
5 898 386 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21216 180
2 5V
-6 -16 8 -8
2 F2
-6 -16 8 -8
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4490 0 0
2
42737.8 1
0
13 Logic Switch~
5 57 33 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21216 0
2 5V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
735 0 0
2
42737.8 0
0
88
1 0 2 0 0 16 0 31 0 0 60 4
206 612
201 612
201 386
463 386
4 2 3 0 0 16 0 36 31 0 0 3
133 315
133 630
206 630
1 3 4 0 0 16 0 36 32 0 0 4
142 269
142 262
167 262
167 240
3 2 5 0 0 16 0 33 36 0 0 2
133 241
133 270
3 3 6 0 0 16 0 34 36 0 0 4
99 241
99 262
124 262
124 269
0 1 7 0 0 16 0 0 32 8 0 3
177 113
176 113
176 195
0 2 8 0 0 16 0 0 32 23 0 3
244 87
158 87
158 195
0 1 7 0 0 16 0 0 33 22 0 3
262 113
142 113
142 196
2 0 8 0 0 16 0 34 0 0 29 2
90 196
90 33
2 0 9 0 0 16 0 33 0 0 11 2
124 196
124 65
2 1 9 0 0 16 0 35 34 0 0 3
158 65
108 65
108 196
1 0 10 0 0 16 0 35 0 0 24 2
194 65
230 65
0 4 11 0 0 16 0 0 10 28 0 3
284 419
436 419
436 453
1 0 12 0 0 16 0 30 0 0 63 3
271 434
271 410
419 410
4 2 13 0 0 16 0 27 30 0 0 2
253 265
253 434
3 2 14 0 0 16 0 31 29 0 0 2
251 621
403 621
3 1 15 0 0 16 0 30 29 0 0 3
262 479
262 603
403 603
3 1 16 0 0 16 0 29 28 0 0 3
449 612
469 612
469 605
1 3 17 0 0 16 0 27 26 0 0 4
262 219
262 166
335 166
335 167
2 3 18 0 0 16 0 27 24 0 0 2
253 220
253 167
3 3 19 0 0 16 0 27 25 0 0 3
244 219
244 167
221 167
1 0 7 0 0 16 0 24 0 0 32 3
262 122
262 113
302 113
2 0 8 0 0 16 0 24 0 0 29 3
244 122
244 87
275 87
1 0 10 0 0 16 0 25 0 0 31 3
230 122
230 65
284 65
2 0 8 0 0 16 0 25 0 0 29 2
212 122
212 33
1 0 7 0 0 16 0 26 0 0 32 2
344 122
344 113
0 2 10 0 0 16 0 0 26 31 0 2
326 64
326 122
3 4 11 0 0 16 0 23 11 0 0 3
284 217
284 453
392 453
2 1 8 0 0 16 0 23 42 0 0 3
275 168
275 33
69 33
1 3 20 0 0 16 0 23 22 0 0 2
293 168
293 173
2 0 10 0 0 16 0 22 0 0 88 3
284 124
284 64
343 64
1 0 7 0 0 16 0 22 0 0 33 3
302 124
302 113
380 113
1 1 7 0 0 16 0 37 1 0 0 4
380 30
380 114
750 114
750 163
2 0 2 0 0 16 0 17 0 0 60 2
732 454
732 386
3 0 21 0 0 16 0 17 0 0 56 2
723 454
723 344
2 0 12 0 0 16 0 16 0 0 63 2
688 454
688 410
3 0 21 0 0 16 0 16 0 0 56 2
679 454
679 344
3 0 22 0 0 16 0 15 0 0 62 2
640 454
640 368
2 0 2 0 0 16 0 15 0 0 60 2
649 454
649 386
3 0 22 0 0 16 0 14 0 0 62 2
597 454
597 368
1 0 12 0 0 16 0 14 0 0 63 2
615 454
615 410
4 0 23 0 0 16 0 17 0 0 45 2
714 454
714 307
4 0 23 0 0 16 0 16 0 0 45 2
670 454
670 307
4 0 23 0 0 16 0 15 0 0 45 2
631 454
631 307
4 1 23 0 0 16 0 14 39 0 0 3
588 454
588 307
884 307
4 0 24 0 0 16 0 13 0 0 61 2
524 454
524 331
3 1 25 0 0 16 0 1 17 0 0 2
741 218
741 454
3 1 26 0 0 16 0 2 16 0 0 3
698 211
697 211
697 454
3 1 27 0 0 16 0 3 15 0 0 2
658 214
658 454
3 2 28 0 0 16 0 4 14 0 0 3
607 211
606 211
606 454
3 3 29 0 0 16 0 6 13 0 0 2
533 212
533 454
3 4 30 0 0 16 0 5 12 0 0 2
482 207
482 454
2 0 21 0 0 16 0 13 0 0 56 2
542 454
542 344
1 0 2 0 0 16 0 13 0 0 60 2
551 454
551 386
3 0 24 0 0 16 0 12 0 0 61 2
491 454
491 331
2 1 21 0 0 16 0 12 40 0 0 3
500 454
500 344
884 344
1 0 12 0 0 16 0 12 0 0 63 2
509 454
509 410
3 0 24 0 0 16 0 10 0 0 61 2
445 453
445 331
0 2 22 0 0 16 0 0 10 62 0 3
455 368
454 368
454 453
1 1 2 0 0 16 0 10 41 0 0 3
463 453
463 386
884 386
2 3 24 0 0 16 0 7 11 0 0 3
832 331
401 331
401 453
2 2 22 0 0 16 0 11 8 0 0 3
410 453
410 368
832 368
2 1 12 0 0 16 0 9 11 0 0 3
832 410
419 410
419 453
5 2 31 0 0 16 0 20 19 0 0 3
470 563
544 563
544 576
5 1 32 0 0 16 0 21 19 0 0 3
667 569
562 569
562 576
1 5 33 0 0 16 0 21 17 0 0 4
680 519
680 516
728 516
728 499
2 5 34 0 0 16 0 21 16 0 0 4
671 519
671 506
684 506
684 499
3 5 35 0 0 16 0 21 15 0 0 4
662 519
662 506
645 506
645 499
4 5 36 0 0 16 0 21 14 0 0 4
653 519
653 515
602 515
602 499
1 5 37 0 0 16 0 20 13 0 0 4
483 513
483 503
538 503
538 499
2 5 38 0 0 16 0 20 12 0 0 3
474 513
474 499
496 499
3 5 39 0 0 16 0 20 10 0 0 3
465 513
465 498
450 498
4 5 40 0 0 16 0 20 11 0 0 5
456 513
456 508
437 508
437 498
406 498
3 1 41 0 0 16 0 19 18 0 0 4
553 622
553 629
497 629
497 605
2 0 10 0 0 16 0 2 0 0 88 2
689 162
689 64
0 1 2 0 0 16 0 0 9 60 0 3
874 386
874 410
868 410
0 1 21 0 0 16 0 0 8 56 0 3
873 344
873 368
868 368
0 1 23 0 0 16 0 0 7 45 0 3
873 307
873 331
868 331
1 0 7 0 0 16 0 2 0 0 33 2
707 162
707 114
1 0 7 0 0 16 0 3 0 0 33 2
667 162
667 114
1 0 7 0 0 16 0 4 0 0 33 2
616 165
616 114
1 0 7 0 0 16 0 6 0 0 33 2
542 161
542 114
1 0 7 0 0 16 0 5 0 0 33 2
491 162
491 114
2 0 10 0 0 16 0 3 0 0 88 3
649 162
650 162
650 64
2 0 10 0 0 16 0 4 0 0 88 2
598 165
598 64
2 0 10 0 0 16 0 6 0 0 88 2
524 161
524 64
2 0 10 0 0 16 0 5 0 0 88 2
473 162
473 64
1 2 10 0 0 16 0 38 1 0 0 4
343 32
343 64
732 64
732 163
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
